library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity InstrMem is
    port(
        A : in std_logic_vector(10 downto 0);
        RD : out std_logic_vector(31 downto 0)
    );
end entity InstrMem;

architecture behavioral of InstrMem is
    type RAM_ARRAY is array (0 to 1023) of std_logic_vector (7 downto 0);
    signal RAM: RAM_ARRAY :=(
        x"00",x"16",x"86",x"93", --addi x13,x13,1  
        x"00",x"56",x"06",x"13", --addi x12,x12,5
        x"00",x"40",x"25",x"03", --lw x10,4(x0)
        x"fe",x"05",x"0e",x"e3", --beq x10,x0,-4
        x"00",x"15",x"85",x"93", --addi x11,x11,1
        x"00",x"c5",x"84",x"63", --beq x11,x12,8
        x"fe",x"00",x"0c",x"e3", --beq x0,x0,-8
        x"00",x"d7",x"0a",x"63", --beq x14,x13,20
        x"00",x"d0",x"20",x"23", --sw x13,0(x0)
        x"40",x"c5",x"85",x"b3", --sub x11,x11,x12
        x"00",x"17",x"07",x"13", --addi x14,x14,1
        x"fe",x"00",x"02",x"e3", --beq x0,x0,-28
        x"00",x"00",x"00",x"00", 
        x"00",x"00",x"20",x"23", --sw x0,0(x0)
        x"40",x"c5",x"85",x"b3", --sub x11,x11,x12
        x"40",x"d7",x"07",x"33", --sub x14,x14,x13
        x"fc",x"00",x"04",x"e3", --beq x0,x0,-56
        x"00",x"00",x"00",x"00", 
        x"00",x"00",x"00",x"00", 
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00"
        ); 
begin
    RD <= RAM(to_integer(signed(A))) & RAM(to_integer(signed(A))+1) & RAM(to_integer(signed(A))+2) & RAM(to_integer(signed(A))+3);
end architecture behavioral;
