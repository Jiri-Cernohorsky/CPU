library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity IOControler is
    port(
        clk : in std_logic;
        rst : in std_logic
    );
end entity IOControler;

architecture behavioral of IOControler is
            
begin

end architecture behavioral;
