library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity InstrMem is
    port(
        A : in std_logic_vector(10 downto 0);
        RD : out std_logic_vector(31 downto 0)
    );
end entity InstrMem;

architecture behavioral of InstrMem is
    type RAM_ARRAY is array (0 to 1023) of std_logic_vector (7 downto 0);
    signal RAM: RAM_ARRAY :=(
        x"40",x"00",x"04",x"93",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"10",x"80",x"93",
        x"00",x"14",x"a0",x"23",
        x"00",x"14",x"a6",x"23",
        x"00",x"13",x"03",x"13",
        x"ff",x"df",x"f0",x"6f",

        x"00",x"10",x"20",x"23",
        x"00",x"20",x"22",x"23",
        x"00",x"30",x"24",x"23",
        x"00",x"40",x"26",x"23",
        x"00",x"50",x"28",x"23",
        x"00",x"60",x"2a",x"23",
        x"00",x"70",x"2c",x"23",
        x"00",x"80",x"2e",x"23",
        x"02",x"90",x"20",x"23",
        x"02",x"a0",x"22",x"23",
        x"02",x"b0",x"24",x"23",
        x"02",x"c0",x"26",x"23",
        x"02",x"d0",x"28",x"23",
        x"02",x"e0",x"2a",x"23",
        x"02",x"f0",x"2c",x"23",
        x"03",x"00",x"2e",x"23",
        x"05",x"10",x"20",x"23",
        x"05",x"20",x"22",x"23",
        x"05",x"30",x"24",x"23",
        x"05",x"40",x"26",x"23",
        x"05",x"50",x"28",x"23",
        x"05",x"60",x"2a",x"23",
        x"05",x"70",x"2c",x"23",
        x"05",x"80",x"2e",x"23",
        x"07",x"90",x"20",x"23",
        x"07",x"a0",x"22",x"23",
        x"07",x"b0",x"24",x"23",
        x"07",x"c0",x"26",x"23",
        x"07",x"d0",x"28",x"23",
        x"07",x"e0",x"2a",x"23",
        x"07",x"f0",x"2c",x"23",
        x"40",x"00",x"04",x"93",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"94",x"84",x"b3",
        x"00",x"84",x"a3",x"03",
        x"00",x"10",x"00",x"93",
        x"00",x"20",x"01",x"13",
        x"00",x"23",x"22",x"33",
        x"00",x"02",x"06",x"63",
        x"00",x"23",x"03",x"33",
        x"00",x"64",x"a4",x"23",
        x"00",x"44",x"a2",x"83",
        x"00",x"12",x"a2",x"33",
        x"00",x"12",x"06",x"63",
        x"00",x"22",x"82",x"b3",
        x"00",x"80",x"00",x"6f",
        x"40",x"22",x"82",x"b3",
        x"00",x"54",x"a2",x"23",
        x"00",x"14",x"a8",x"23",
        x"00",x"00",x"20",x"83",
        x"00",x"40",x"21",x"03",
        x"00",x"80",x"21",x"83",
        x"00",x"c0",x"22",x"03",
        x"01",x"00",x"22",x"83",
        x"01",x"40",x"23",x"03",
        x"01",x"80",x"23",x"83",
        x"01",x"c0",x"24",x"03",
        x"02",x"00",x"24",x"83",
        x"02",x"40",x"25",x"03",
        x"02",x"80",x"25",x"83",
        x"02",x"c0",x"26",x"03",
        x"03",x"00",x"26",x"83",
        x"03",x"40",x"27",x"03",
        x"03",x"80",x"27",x"83",
        x"03",x"c0",x"28",x"03",
        x"04",x"00",x"28",x"83",
        x"04",x"40",x"29",x"03",
        x"04",x"80",x"29",x"83",
        x"04",x"c0",x"2a",x"03",
        x"05",x"00",x"2a",x"83",
        x"05",x"40",x"2b",x"03",
        x"05",x"80",x"2b",x"83",
        x"05",x"c0",x"2c",x"03",
        x"06",x"00",x"2c",x"83",
        x"06",x"40",x"2d",x"03",
        x"06",x"80",x"2d",x"83",
        x"06",x"c0",x"2e",x"03",
        x"07",x"00",x"2e",x"83",
        x"07",x"40",x"2f",x"03",
        x"07",x"80",x"2f",x"83",
        x"30",x"20",x"00",x"73",
        x"00",x"00",x"00",x"00", 
        x"00",x"00",x"00",x"00", 
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00",
        x"00",x"00",x"00",x"00"
        ); 
begin
    RD <= RAM(to_integer(signed(A))) & RAM(to_integer(signed(A))+1) & RAM(to_integer(signed(A))+2) & RAM(to_integer(signed(A))+3);
end architecture behavioral;
